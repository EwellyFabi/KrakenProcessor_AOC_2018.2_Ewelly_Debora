library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity KrakenProcessor is

port( 
	clock : in std_logic
 );
    
end KrakenProcessor;

architecture kraken of KrakenProcessor is
begin



end kraken;